`include "mux.v"

`include "prj_definition.v"
module MUX32_32x1_TB;

  reg[`DATA_INDEX_LIMIT:0] I0, I1, I2, I3, I4, I5, I6, I7,
                           I8, I9, I10, I11, I12, I13, I14, I15,
                           I16, I17, I18, I19, I20, I21, I22, I23,
                           I24, I25, I26, I27, I28, I29, I30, I31;
  reg[4:0] S;
  wire[`DATA_INDEX_LIMIT:0] Y;
  MUX32_32x1 MUX32_32x1_INST(Y, I0, I1, I2, I3, I4, I5, I6, I7,
                                I8, I9, I10, I11, I12, I13, I14, I15,
                                I16, I17, I18, I19, I20, I21, I22, I23,
                                I24, I25, I26, I27, I28, I29, I30, I31, S);

  initial begin
    $dumpfile("tb.vcd");
    $dumpvars(0, MUX32_32x1_TB);
    S='b00000;I0='h00000000;I1='h00000000;I2='h00000000;I3='h00000000;I4='h00000000;I5='h00000000;I6='h00000000;I7='h00000000;
            I8='h88888888;I9='h99999999;I10='haaaa1010;I11='hbbbb1111;I12='hcccc1212;I13='hdddd1313;I14='heeee1414;I15='hffff1515;
            I16='h16161616;I17='h17171717;I18='h18181818;I19='h19191919;I20='h20202020;I21='h21212121;I22='h22222222;I23='h23232323;
            I24='h24242424;I25='h25252525;I26='h26262626;I27='h27272727;I28='h28282828;I29='h29292929;I30='h30303030;I31='h31313131;
    #5 S='b00000;I0='h00012340;I1='habc21000;I2='h00033300;I3='h00aadd00;I4='h44444444;I5='h55555555;I6='h66666666;I7='h77777777;
    #5 S='b00001;I0='h22330000;I1='hffffffff;I2='h9999ffdd;I3='h00000001;I4='h44444444;I5='h55555555;I6='h66666666;I7='h77777777;
    #5 S='b00010;I0='h00001230;I1='h02220000;I2='h0000ade0;I3='h00000000;I4='h44444444;I5='h55555555;I6='h66666666;I7='h77777777;
    #5 S='b00011;I0='h09090901;I1='h0000efd1;I2='h94588255;I3='hacdefb00;I4='h44444444;I5='h55555555;I6='h66666666;I7='h77777777;
    #5 S='b00100;I0='h00000000;I1='h00000001;I2='h00000002;I3='h00000003;I4='h44444444;I5='h55555555;I6='h66666666;I7='h77777777;
    #5 S='b00101;I0='h00000000;I1='h00000001;I2='h00000002;I3='h00000003;I4='h44444444;I5='h55555555;I6='h66666666;I7='h77777777;
    #5 S='b00110;I0='h00000000;I1='h00000001;I2='h00000002;I3='h00000003;I4='h44444444;I5='h55555555;I6='h66666666;I7='h77777777;
    #5 S='b00111;I0='h00000000;I1='h00000001;I2='h00000002;I3='h00000003;I4='h44444444;I5='h55555555;I6='h66666666;I7='h77777777;
    #5 S='b01000;
    #5 S='b01001;
    #5 S='b01010;
    #5 S='b01011;
    #5 S='b01100;
    #5 S='b01101;
    #5 S='b01110;
    #5 S='b01111;
    #5 S='b10000;
    #5 S='b10001;
    #5 S='b10010;
    #5 S='b10011;
    #5 S='b10100;
    #5 S='b10101;
    #5 S='b10110;
    #5 S='b10111;
    #5 S='b11000;
    #5 S='b11001;
    #5 S='b11010;
    #5 S='b11011;
    #5 S='b11100;
    #5 S='b11101;
    #5 S='b11110;
    #5 S='b11111;
    #5
    $finish;
  end

endmodule
