`include "mux.v"

`include "prj_definition.v"
module MUX1_32x1_TB;

  reg I0, I1, I2, I3, I4, I5, I6, I7,
      I8, I9, I10, I11, I12, I13, I14, I15,
      I16, I17, I18, I19, I20, I21, I22, I23,
      I24, I25, I26, I27, I28, I29, I30, I31;
  reg [4:0]S;
  wire Y;
  MUX1_32x1 MUX1_32x1_INST(Y, I0, I1, I2, I3, I4, I5, I6, I7,
                              I8, I9, I10, I11, I12, I13, I14, I15,
                              I16, I17, I18, I19, I20, I21, I22, I23,
                              I24, I25, I26, I27, I28, I29, I30, I31, S);

  initial begin
    $dumpfile("tb.vcd");
    $dumpvars(0, MUX1_32x1_TB);
    S='b00000;I0=1;I1=0;I2=1;I3=0;I4=1;I5=0;I6=1;I7=0;I8=1;I9=0;I10=1;I11=0;I12=1;I13=0;I14=1;I15=0;
             I16=1;I17=0;I18=1;I19=0;I20=1;I21=0;I22=1;I23=0;I24=1;I25=0;I26=1;I27=0;I28=1;I29=0;I30=1;I31=0;
    #5 S='b00000;
    #5 S='b00001;
    #5 S='b00010;
    #5 S='b00011;
    #5 S='b00100;
    #5 S='b00101;
    #5 S='b00110;
    #5 S='b00111;
    #5 S='b01000;
    #5 S='b01001;
    #5 S='b01010;
    #5 S='b01011;
    #5 S='b01100;
    #5 S='b01101;
    #5 S='b01110;
    #5 S='b01111;
    #5 S='b10000;
    #5 S='b10001;
    #5 S='b10010;
    #5 S='b10011;
    #5 S='b10100;
    #5 S='b10101;
    #5 S='b10110;
    #5 S='b10111;
    #5 S='b11000;
    #5 S='b11001;
    #5 S='b11010;
    #5 S='b11011;
    #5 S='b11100;
    #5 S='b11101;
    #5 S='b11110;
    #5 S='b11111;
    #5
    $finish;
  end

endmodule
